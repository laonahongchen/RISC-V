module if (
    input wire[`InstAddrBus] pc,
    input wire[`InstBus] inst,
    output reg pc_o,
    output reg inst_o,
    output reg stall_req_o
);

endmodule // if
